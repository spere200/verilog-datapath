`include "SignExtend.v"
`include "Control.v"
`include "ALUControl.v"
`include "ALU.v"
`include "Adder.v"
`include "Incrementer.v"
`include "PCSelector.v"
`include "Shifter.v"
`include "Mux3to1.v"

module Datapath;
	////////////////////
	////clock signal////
	////////////////////
	reg clock;
	
	initial begin
		clock = 0;
	end
	
	always begin
		#20 clock = ~clock;
	end
	
	////////////////////
	//end clock signal//
	////////////////////
	
	/////////////////////////////////////////////////////////////////////////////////////
	////////////////////////////BEGIN DECLARATION BLOCK//////////////////////////////////
	/////////////////////////////////////////////////////////////////////////////////////
	
	//single registers
	reg [63:0] PC;
	
	reg HazardBit;
	
	//pipeline registers
	reg [95 :0]	IFID;
	reg [291:0]	IDEX; //IDEX was expanded to store Reg1 and Reg2 (source reg. addresses)
	reg [204:0]	EXMEM;
	reg [135:0]	MEMWB; //increased to store written data
	
	//control signal wires
	wire [3:0] ALUctl;
	wire [1:0] ALUOp;
	wire Reg2Loc, Uncondbranch, nzBranch, zBranch, MemRead, MemtoReg, MemWrite, 
		 ALUSrc, RegWrite;
	wire PCSrc; //not generated by the control, determines source of PC
	
	//data transfer wires
	wire [63:0] ALUInA, ALUInB, ALUOut, FwdALUInA, FwdALUInB; 
	reg  [1:0 ] FwdASelector, FwdBSelector;
	wire [63:0] ExtendedOffset; //sign extended offset
	wire [63:0] IncrementedPC, BranchPC, PCValue; //wires used for calculating next PC
	wire [63:0] RWriteData; //data being written to the target register
	wire [63:0] PCAdderInputB; //ExtendedOffset shifted to the left twice
	wire [63:0] MemWriteData; //data being written to memory
	wire [63:0] Reg2Data, Reg1Data;
	wire [4:0 ]  Reg2, Reg1; //address of source registers
	wire Zero; //zero signal of the ALU
	
	//declaring register file, instruction memory, and data memory
	reg [63:0] RF[31:0]; //32 registers each 64 bits long
	reg [7:0] MDR[8191:0]; //8192 bytes (1024 doublewords)
	reg [7:0] MIR[4095:0]; //4096 bytes (1024 words)
	
	//integer i;
	
	//Begin loading Instruction Memory and Data Memory
	initial begin 
		$readmemh("IM_Extra_Bytes.txt", MIR);
		$readmemh("DM_Bytes.txt", MDR);
		
		//initialize pipeline registers
		IFID <= 0;
		IDEX <= 0;
		EXMEM <= 0;
		MEMWB <= 0;
		
		PC <= 0;
		HazardBit <= 0;
	end
	//End loading Instruction Memory and Data Memory
	
	
	/////////////////////////////////////////////////////////////////////////////////////
	//////////////////////////////END DECLARATION BLOCK//////////////////////////////////
	/////////////////////////////////////////////////////////////////////////////////////
	
	/////////////////////////////////////////////////////////////////////////////////////
	///////////////////////////BEGIN COMBINATIONAL BLOCK/////////////////////////////////
	/////////////////////////////////////////////////////////////////////////////////////
	
	//wires value assignment w/ multiplexers
	assign Reg1 = IFID[9:5];
	assign Reg2 = IFID[28] ? IFID[4:0] : IFID[20:16]; //Reg2Loc replaced by Instruction[28]
	assign Reg1Data = RF[Reg1];
	assign Reg2Data = RF[Reg2];
	assign ALUInA = IDEX[207:144];
	assign ALUInB = IDEX[279] ? IDEX[79:16] : IDEX[143:80]; //ALUSrc replaced by IDEX[279]
	assign PCSrc = (EXMEM[204] || (EXMEM[203] && EXMEM[133]) || (EXMEM[202] && ~EXMEM[133])) ? 1 : 0;
	
	//shift ExtendedOffset 2 to the left and save it in PCAdderInputB
	Shifter shiftOffset(IDEX[79:16], PCAdderInputB);
	
	//control signal generation
	Control controller(IFID[31:21], Reg2Loc, Uncondbranch, nzBranch, zBranch, 
							  MemRead, MemtoReg, ALUOp, MemWrite, ALUSrc, RegWrite);
		
	//ALU operations
	SignExtend extender(IFID[31:0], ExtendedOffset); //extend offset field
	ALUControl ALUC(IDEX[281:280], IDEX[15:5], ALUctl);
	ALU alu(ALUctl, FwdALUInA, FwdALUInB, ALUOut, Zero);

	//PC calculation
	Incrementer incrPC(PC, IncrementedPC); //calculate incremented PC
	Adder branPC(IDEX[271:208], PCAdderInputB, BranchPC); //calculate branched PC
	
	//setting PC
	PCSelector pcval(PCSrc, EXMEM[197:134], IncrementedPC, PCValue);
	
	/////////////////////////////////////////////////////////////////////////////////////
	////////////////////////////END COMBINATIONAL BLOCK//////////////////////////////////
	/////////////////////////////////////////////////////////////////////////////////////
	
	/////////////////////////////////////////////////////////////////////////////////////
	/////////////////////////////////BEGIN FORWARDING////////////////////////////////////
	/////////////////////////////////////////////////////////////////////////////////////
	
	//3-to-1 multiplexers to select the correct ALU inputs (normal, EXMEM, or MEMWB)
	Mux3to1 aForward(FwdASelector, ALUInA, MEMWB[68:5], EXMEM[132:69], MEMWB[132:69], FwdALUInA);
	Mux3to1 bForward(FwdBSelector, ALUInB, MEMWB[68:5], EXMEM[132:69], MEMWB[132:69], FwdALUInB);
	
	always @(PC, IDEX, EXMEM, MEMWB) begin
		
		//Setting selector for A forwarding
		if(IDEX[15:5] != 1704) begin
			if( (EXMEM[4:0] != 31) && (EXMEM[4:0] == IDEX[291:287]) && (EXMEM[198]) ) begin
				FwdASelector <= 2;
			end
			else if( (MEMWB[4:0] != 31) && (MEMWB[4:0] == IDEX[291:287]) && (MEMWB[133]) && (MEMWB[135]) ) begin
				FwdASelector <= 3;
			end
			else if( (MEMWB[4:0] != 31) && (MEMWB[4:0] == IDEX[291:287]) && (MEMWB[133]) && ~(MEMWB[135]) ) begin
				FwdASelector <= 1;
			end
			else begin FwdASelector = 0; end
			
			//Setting selector for B forwarding
			if(~IDEX[274]) begin //if it's not a STUR
				if( (EXMEM[4:0] != 31) && (EXMEM[4:0] == IDEX[286:282]) && (EXMEM[198]) ) begin
					FwdBSelector <= 2;
				end
				
				else if( (MEMWB[4:0] != 31) && (MEMWB[4:0] == IDEX[286:282]) && (MEMWB[133]) && (MEMWB[135]) ) begin
					FwdBSelector <= 3;
				end
				
				else if( (MEMWB[4:0] != 31) && (MEMWB[4:0] == IDEX[286:282]) && (MEMWB[133]) && ~(MEMWB[135]) ) begin
					FwdBSelector <= 1;
				end
				
				else begin
					FwdBSelector <= 0; 	
				end
			end
			
			//for STUR, forwarding the second value needs to be done differently, since STUR uses the forwarded
			//value as-is, it doesn't use it for ALU operations. Forwarding is done directly
			else begin
				if( (EXMEM[4:0] != 31) && (EXMEM[4:0] == IDEX[4:0]) && (EXMEM[198]) ) begin
					FwdBSelector <= 0;
					IDEX[143:80] <= EXMEM[132:69];
				end
				
				else if( (MEMWB[4:0] != 31) && (MEMWB[4:0] == IDEX[4:0]) && (MEMWB[133]) && (MEMWB[135]) ) begin
					FwdBSelector <= 0;
					IDEX[143:80] <= MEMWB[132:69];
				end
				
				else if( (MEMWB[4:0] != 31) && (MEMWB[4:0] == IDEX[4:0]) && (MEMWB[133]) && ~(MEMWB[135]) ) begin
					FwdBSelector <= 0;
					IDEX[143:80] <= MEMWB[68:5];
				end
				
				else begin
					FwdBSelector <= 0;
				end
			end
		end
	end
	
	//Data Hazard check, only used for read after LDUR to
	//delay the instruction by inserting a bubble
	always @(PC, IFID, IDEX) begin
		if(IDEX[275]) begin
			if(IDEX[4:0] == Reg1) begin
				HazardBit <= 1;
				IFID[31:0] <= 32'hD503201F;
			end
			
			//only check Reg2 if Reg2Loc is 0 (R-Type)
			if((MemtoReg == 0) && (IFID[28] == 0)) begin
				HazardBit <= 1;
				IFID[31:0] <= 32'hD503201F;
			end
		end
	end
	
	/////////////////////////////////////////////////////////////////////////////////////
	/////////////////////////////////END FORWARDING//////////////////////////////////////
	/////////////////////////////////////////////////////////////////////////////////////
		
	/////////////////////////////////////////////////////////////////////////////////////
	////////////////////////////BEGIN SEQUENTIAL BLOCK///////////////////////////////////
	/////////////////////////////////////////////////////////////////////////////////////
	
	//if instruction is HALT dump output file and finish
	always @(IFID) begin
		if(IFID[31:21] == {11{1'b1}}) 
			begin 
				//output the data memory to a new file and end simulation
				$writememh("DM_Final_Bytes.txt", MDR);
				$finish;
			end
	end
	
	always @(MEMWB, EXMEM) begin
		//writing to memory or register on clock edge
		if (MEMWB[133]) begin
			if(MEMWB[134]) begin RF[MEMWB[4:0]] <= MEMWB[132:69]; end
			else		   begin RF[MEMWB[4:0]] <= MEMWB[68 : 5]; end
		end
		
		if(EXMEM[200]) begin
			MDR[EXMEM[132: 69]    ] <= EXMEM[12: 5];
			MDR[EXMEM[132: 69] + 1] <= EXMEM[20:13];
			MDR[EXMEM[132: 69] + 2] <= EXMEM[28:21];
			MDR[EXMEM[132: 69] + 3] <= EXMEM[36:29];
			MDR[EXMEM[132: 69] + 4] <= EXMEM[44:37];
			MDR[EXMEM[132: 69] + 5] <= EXMEM[52:45];
			MDR[EXMEM[132: 69] + 6] <= EXMEM[60:53];
			MDR[EXMEM[132: 69] + 7] <= EXMEM[68:61];
		end
	end
	
	
	always @(PC) begin
		#1 $display("PC: %3d  Instr: %8h  A: %3d  B: %3d  Out: %3d  X7: %3d", IFID[95:32], IFID[31:0], $signed(FwdALUInA), $signed(FwdALUInB), $signed(ALUOut), $signed(RF[7]));
	end
	
	//clock dependent logic
	//each clock cycle a new instruction is fetched
	//and instructions in the pipeline move up
	always @(posedge clock) begin
		//Ground XZR
		RF[31] = 0;
		
		//HAZARD CHECKING CODE
		if(HazardBit == 0) begin
			PC <= PCValue;
		end
		else begin
			HazardBit <= 0;
			PC <= PC;
		end
		
		//IFID steps
		IFID[95:32] <= PC;
		IFID[ 7: 0] <= MIR[PC    ];
		IFID[15: 8] <= MIR[PC + 1];
		IFID[23:16] <= MIR[PC + 2];
		IFID[31:24] <= MIR[PC + 3];
		
		//IDEX steps w/ hazard checking
		if(HazardBit) begin
			IDEX[281:280] <= 0;
			IDEX[279	] <= 0;
			IDEX[278	] <= 0;
			IDEX[277	] <= 0;
			IDEX[276	] <= 0;
			IDEX[275	] <= 0;
			IDEX[274	] <= 0;
			IDEX[273	] <= 0;
			IDEX[272	] <= 0;
		end
		
		else begin
			IDEX[281:280] <= ALUOp;			//storing necessary control signals
			IDEX[279	] <= ALUSrc;
			IDEX[278	] <= Uncondbranch;
			IDEX[277	] <= zBranch;
			IDEX[276	] <= nzBranch;
			IDEX[275	] <= MemRead;
			IDEX[274	] <= MemWrite;
			IDEX[273	] <= MemtoReg;
			IDEX[272	] <= RegWrite;
		end
		//end hazard correction in IDEX
		
		IDEX[271:208] <= IFID[95:32];
		IDEX[207:144] <= Reg1Data;
		IDEX[143: 80] <= Reg2Data;
		IDEX[79 : 16] <= ExtendedOffset;
		IDEX[15 :  5] <= IFID[31:21];
		IDEX[4  :  0] <= IFID[4:0]; //store Rt/Rd
		IDEX[291:287] <= Reg1; //store Rm
		IDEX[286:282] <= Reg2; //store Rn
		
		//EXMEM steps
		EXMEM[204	] <= IDEX[278];		//storing necessary control signals
		EXMEM[203	] <= IDEX[277];
		EXMEM[202	] <= IDEX[276];
		EXMEM[201	] <= IDEX[275];
		EXMEM[200	] <= IDEX[274];
		EXMEM[199	] <= IDEX[273];
		EXMEM[198	] <= IDEX[272];
		
		EXMEM[197:134] <= BranchPC;
		EXMEM[133    ] <= Zero;
		EXMEM[132: 69] <= ALUOut;
		EXMEM[68 :  5] <= IDEX[143:80];
		EXMEM[4  :  0] <= IDEX[4:0];
		
		//MEMWB steps
		MEMWB[134] <= EXMEM[199];		//storing necessary control signals
		MEMWB[133] <= EXMEM[198];
		
		MEMWB[132:125] <= MDR[EXMEM[132:69] + 7];	//array read from memory
		MEMWB[124:117] <= MDR[EXMEM[132:69] + 6];
		MEMWB[116:109] <= MDR[EXMEM[132:69] + 5];
		MEMWB[108:101] <= MDR[EXMEM[132:69] + 4];
		MEMWB[100: 93] <= MDR[EXMEM[132:69] + 3];
		MEMWB[92 : 85] <= MDR[EXMEM[132:69] + 2];
		MEMWB[84 : 77] <= MDR[EXMEM[132:69] + 1];
		MEMWB[76 : 69] <= MDR[EXMEM[132:69]    ];
		
		MEMWB[68 :  5] <= EXMEM[132:69];
		
		MEMWB[4  :  0] <= EXMEM[4:0];
		
		MEMWB[135    ] <= EXMEM[201];
	end
	/////////////////////////////////////////////////////////////////////////////////////
	/////////////////////////////END SEQUENTIAL BLOCK////////////////////////////////////
	/////////////////////////////////////////////////////////////////////////////////////
endmodule